//module tb_fir;
//
//	logic clk_05;
//	logic rst;
//	logic CLOCK_50;
//	logic [0:0]SW;
////	logic signed [15:0] in;
////	logic input_ready;
//	logic signed [15:0] out;
//	logic output_ready;
//	
//	int count = 0;
//	
//
//	FIR CUT (.*);
//	
//	initial
//		begin
//			SW=1;
//
//			clk_05=0;
//			rst = 1;
//		end
//		
//	always
//		begin
//			#20ns clk_05=~clk_05;
//		end
//		
//	always 
//		begin
//			
//		#100ns;
//		
//		SW=1;
//		
//		#100ns;
//		
//		SW=1;
//		
//		end	
//
//endmodule
